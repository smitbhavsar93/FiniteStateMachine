library verilog;
use verilog.vl_types.all;
entity fsm_vlg_vec_tst is
end fsm_vlg_vec_tst;
